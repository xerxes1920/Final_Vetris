module rx(
	input clk,
	input rst,
	//input iocs,
    //input iorw,
    input rxd,
    input rate_en,
	input [1:0] ioaddr,
    input [7:0] rx_ack,

    output reg rda,
    output reg [7:0] rx2bus
    ); 

    parameter IO_XFER=2'b00, REG_RD=2'b01, LD_DIV_LO=2'b10, LD_DIV_HI=2'b11;
	parameter WAIT=3'b000, START_L=3'b001, DATA=3'b010, STOP=3'b100; 

    reg [2:0] state;
	reg [2:0] nxt_state;    

	reg shift;  		//if need to shift bit
	reg rst_per; 		//if need to reset period 
	reg clr_bit_cnt;	//clear bit counter
	reg inc_bit_cnt;	//inc bit counter
    reg set_rdy;		//ready!
    reg clr_rdy;
    reg [2:0] bit_cnt;

    //state register
	always @ (posedge clk or negedge rst) begin
		if(!rst)
			state = WAIT;
		else
			state = nxt_state;
	end
		

	//RX shift register
	always @ (posedge clk)
		if (!rst)
	    rx2bus <= 8'h00;
	  else if (shift)
	    rx2bus <= {rxd,rx2bus[7:1]};
	
	
	//bit counter 
	always @ (posedge clk)
	  if (clr_bit_cnt)
	    bit_cnt <= 3'b000;
	  else if (inc_bit_cnt)
	    bit_cnt <= bit_cnt + 3'b001;

	//rdy flop //
	always @ (posedge clk)
		if (!rst)
	    rda <= 1'b0;
	  else if (set_rdy)
	    rda <= 1'b1;
	  else if (clr_rdy)
	    rda <= 1'b0;

    //RX SM
	always@(*) begin
		//Set defaults
		shift = 1'b0;
		rst_per = 1'b0;
		clr_bit_cnt = 1'b0;
		inc_bit_cnt = 1'b0;
		set_rdy = 1'b0;
		clr_rdy = 1'b0;
		nxt_state = state;
		
		case (state)
		  WAIT: begin
		    clr_rdy = 1'b1;
            if(ioaddr == IO_XFER) begin
                //clr_rdy = 1'b1;
                clr_bit_cnt = 1'b1;
                nxt_state = START_L;
            end
          end
	 	  START_L : begin //Looking for the start bit
		    if ((rxd == 1'b0) && rate_en) begin
			  nxt_state = DATA;
			end /*else if(RX == 1'b1) begin
				nxt_state = IDLE;
		  end*/ 
		  //shrink it for size
		  end
		  DATA : begin //recieving
		   if (rate_en) begin
				inc_bit_cnt = 1'b1;
				shift = 1'b1;
				nxt_state = (&bit_cnt)?STOP:DATA;
			 end
		  end
          default: begin //same as stop, wait for a period for the stop bit
          	if (rate_en) begin
			  nxt_state = WAIT;
              set_rdy = 1'b1;
          	end
		  end
		endcase
	end
endmodule
