module MP2Graphics(
    clk,
    rst,
    oData,
    dVal
);

input logic clk, rst, dVal;
input logic [35:0] oData;

output logic dVal;



endmodule
